library verilog;
use verilog.vl_types.all;
entity testall is
end testall;
