library verilog;
use verilog.vl_types.all;
entity test_fsm is
end test_fsm;
