library verilog;
use verilog.vl_types.all;
entity test_regs is
end test_regs;
