module pc(clk,npc,reset,pcout);
  input clk,reset;
  input [31:0] npc;
  output [31:0] pcout;
  reg [31:0] pcout;
  
  
  always @(posedge clk,posedge reset)
  begin
    if(reset)//reset=1 ??
      pcout=32'h0000_3000;
    else
      pcout<=npc;
  end
endmodule