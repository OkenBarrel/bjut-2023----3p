library verilog;
use verilog.vl_types.all;
entity bgetest is
end bgetest;
